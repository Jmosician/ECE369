module TopLevel(Clk, Rst, PCValue,WriteData);
    input Clk,Rst;
    output [31:0] PCValue;
    output [31:0] WriteData;












endmodule